/* ds */ 
